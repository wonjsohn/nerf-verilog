module waveform_from_lut(clk, reset, value);
input wire          clk;
input wire          reset;
output reg [31:0]   value;

// *** Declarations
reg [9:0]    index;


	always @ (posedge clk or posedge reset) begin
        if (reset) begin
            index <= 10'd0;
            value <= 32'h3f4ccccd;
        end
        else begin // not reset
            if (index == 10'd1023) begin
                index <= 10'd0;
            end
            else begin // index < maxlength
                index <= index + 10'd1;
            end
            case (index)                
                10'd0  : value <= 32'h3f4ccccd;
                10'd1  : value <= 32'h3f4ccd0c;
                10'd2  : value <= 32'h3f4ccdca;
                10'd3  : value <= 32'h3f4ccf06;
                10'd4  : value <= 32'h3f4cd0c1;
                10'd5  : value <= 32'h3f4cd2fb;
                10'd6  : value <= 32'h3f4cd5b3;
                10'd7  : value <= 32'h3f4cd8e9;
                10'd8  : value <= 32'h3f4cdc9e;
                10'd9  : value <= 32'h3f4ce0d2;
                10'd10  : value <= 32'h3f4ce584;
                10'd11  : value <= 32'h3f4ceab4;
                10'd12  : value <= 32'h3f4cf062;
                10'd13  : value <= 32'h3f4cf68f;
                10'd14  : value <= 32'h3f4cfd3a;
                10'd15  : value <= 32'h3f4d0463;
                10'd16  : value <= 32'h3f4d0c0a;
                10'd17  : value <= 32'h3f4d142f;
                10'd18  : value <= 32'h3f4d1cd2;
                10'd19  : value <= 32'h3f4d25f2;
                10'd20  : value <= 32'h3f4d2f91;
                10'd21  : value <= 32'h3f4d39ad;
                10'd22  : value <= 32'h3f4d4446;
                10'd23  : value <= 32'h3f4d4f5d;
                10'd24  : value <= 32'h3f4d5af1;
                10'd25  : value <= 32'h3f4d6703;
                10'd26  : value <= 32'h3f4d7391;
                10'd27  : value <= 32'h3f4d809d;
                10'd28  : value <= 32'h3f4d8e25;
                10'd29  : value <= 32'h3f4d9c2a;
                10'd30  : value <= 32'h3f4daaac;
                10'd31  : value <= 32'h3f4db9aa;
                10'd32  : value <= 32'h3f4dc924;
                10'd33  : value <= 32'h3f4dd91b;
                10'd34  : value <= 32'h3f4de98d;
                10'd35  : value <= 32'h3f4dfa7c;
                10'd36  : value <= 32'h3f4e0be6;
                10'd37  : value <= 32'h3f4e1dcb;
                10'd38  : value <= 32'h3f4e302c;
                10'd39  : value <= 32'h3f4e4308;
                10'd40  : value <= 32'h3f4e565f;
                10'd41  : value <= 32'h3f4e6a31;
                10'd42  : value <= 32'h3f4e7e7d;
                10'd43  : value <= 32'h3f4e9344;
                10'd44  : value <= 32'h3f4ea884;
                10'd45  : value <= 32'h3f4ebe3f;
                10'd46  : value <= 32'h3f4ed474;
                10'd47  : value <= 32'h3f4eeb22;
                10'd48  : value <= 32'h3f4f024a;
                10'd49  : value <= 32'h3f4f19ea;
                10'd50  : value <= 32'h3f4f3204;
                10'd51  : value <= 32'h3f4f4a96;
                10'd52  : value <= 32'h3f4f63a1;
                10'd53  : value <= 32'h3f4f7d23;
                10'd54  : value <= 32'h3f4f971e;
                10'd55  : value <= 32'h3f4fb190;
                10'd56  : value <= 32'h3f4fcc7a;
                10'd57  : value <= 32'h3f4fe7db;
                10'd58  : value <= 32'h3f5003b3;
                10'd59  : value <= 32'h3f502002;
                10'd60  : value <= 32'h3f503cc6;
                10'd61  : value <= 32'h3f505a01;
                10'd62  : value <= 32'h3f5077b2;
                10'd63  : value <= 32'h3f5095d8;
                10'd64  : value <= 32'h3f50b474;
                10'd65  : value <= 32'h3f50d384;
                10'd66  : value <= 32'h3f50f309;
                10'd67  : value <= 32'h3f511303;
                10'd68  : value <= 32'h3f513370;
                10'd69  : value <= 32'h3f515451;
                10'd70  : value <= 32'h3f5175a5;
                10'd71  : value <= 32'h3f51976d;
                10'd72  : value <= 32'h3f51b9a7;
                10'd73  : value <= 32'h3f51dc54;
                10'd74  : value <= 32'h3f51ff72;
                10'd75  : value <= 32'h3f522303;
                10'd76  : value <= 32'h3f524705;
                10'd77  : value <= 32'h3f526b77;
                10'd78  : value <= 32'h3f52905b;
                10'd79  : value <= 32'h3f52b5af;
                10'd80  : value <= 32'h3f52db73;
                10'd81  : value <= 32'h3f5301a6;
                10'd82  : value <= 32'h3f532849;
                10'd83  : value <= 32'h3f534f5a;
                10'd84  : value <= 32'h3f5376da;
                10'd85  : value <= 32'h3f539ec8;
                10'd86  : value <= 32'h3f53c724;
                10'd87  : value <= 32'h3f53efed;
                10'd88  : value <= 32'h3f541923;
                10'd89  : value <= 32'h3f5442c6;
                10'd90  : value <= 32'h3f546cd5;
                10'd91  : value <= 32'h3f54974f;
                10'd92  : value <= 32'h3f54c235;
                10'd93  : value <= 32'h3f54ed86;
                10'd94  : value <= 32'h3f551941;
                10'd95  : value <= 32'h3f554566;
                10'd96  : value <= 32'h3f5571f5;
                10'd97  : value <= 32'h3f559eed;
                10'd98  : value <= 32'h3f55cc4e;
                10'd99  : value <= 32'h3f55fa17;
                10'd100  : value <= 32'h3f562848;
                10'd101  : value <= 32'h3f5656e0;
                10'd102  : value <= 32'h3f5685e0;
                10'd103  : value <= 32'h3f56b546;
                10'd104  : value <= 32'h3f56e512;
                10'd105  : value <= 32'h3f571544;
                10'd106  : value <= 32'h3f5745db;
                10'd107  : value <= 32'h3f5776d6;
                10'd108  : value <= 32'h3f57a836;
                10'd109  : value <= 32'h3f57d9fa;
                10'd110  : value <= 32'h3f580c20;
                10'd111  : value <= 32'h3f583eaa;
                10'd112  : value <= 32'h3f587196;
                10'd113  : value <= 32'h3f58a4e4;
                10'd114  : value <= 32'h3f58d892;
                10'd115  : value <= 32'h3f590ca2;
                10'd116  : value <= 32'h3f594112;
                10'd117  : value <= 32'h3f5975e2;
                10'd118  : value <= 32'h3f59ab11;
                10'd119  : value <= 32'h3f59e09f;
                10'd120  : value <= 32'h3f5a168b;
                10'd121  : value <= 32'h3f5a4cd5;
                10'd122  : value <= 32'h3f5a837c;
                10'd123  : value <= 32'h3f5aba80;
                10'd124  : value <= 32'h3f5af1e0;
                10'd125  : value <= 32'h3f5b299b;
                10'd126  : value <= 32'h3f5b61b2;
                10'd127  : value <= 32'h3f5b9a23;
                10'd128  : value <= 32'h3f5bd2ee;
                10'd129  : value <= 32'h3f5c0c12;
                10'd130  : value <= 32'h3f5c458f;
                10'd131  : value <= 32'h3f5c7f65;
                10'd132  : value <= 32'h3f5cb993;
                10'd133  : value <= 32'h3f5cf417;
                10'd134  : value <= 32'h3f5d2ef3;
                10'd135  : value <= 32'h3f5d6a24;
                10'd136  : value <= 32'h3f5da5ab;
                10'd137  : value <= 32'h3f5de187;
                10'd138  : value <= 32'h3f5e1db7;
                10'd139  : value <= 32'h3f5e5a3b;
                10'd140  : value <= 32'h3f5e9712;
                10'd141  : value <= 32'h3f5ed43c;
                10'd142  : value <= 32'h3f5f11b7;
                10'd143  : value <= 32'h3f5f4f84;
                10'd144  : value <= 32'h3f5f8da2;
                10'd145  : value <= 32'h3f5fcc11;
                10'd146  : value <= 32'h3f600ace;
                10'd147  : value <= 32'h3f6049db;
                10'd148  : value <= 32'h3f608936;
                10'd149  : value <= 32'h3f60c8df;
                10'd150  : value <= 32'h3f6108d5;
                10'd151  : value <= 32'h3f614918;
                10'd152  : value <= 32'h3f6189a7;
                10'd153  : value <= 32'h3f61ca81;
                10'd154  : value <= 32'h3f620ba5;
                10'd155  : value <= 32'h3f624d14;
                10'd156  : value <= 32'h3f628ecc;
                10'd157  : value <= 32'h3f62d0cd;
                10'd158  : value <= 32'h3f631316;
                10'd159  : value <= 32'h3f6355a7;
                10'd160  : value <= 32'h3f63987e;
                10'd161  : value <= 32'h3f63db9c;
                10'd162  : value <= 32'h3f641eff;
                10'd163  : value <= 32'h3f6462a7;
                10'd164  : value <= 32'h3f64a693;
                10'd165  : value <= 32'h3f64eac3;
                10'd166  : value <= 32'h3f652f36;
                10'd167  : value <= 32'h3f6573ec;
                10'd168  : value <= 32'h3f65b8e2;
                10'd169  : value <= 32'h3f65fe1a;
                10'd170  : value <= 32'h3f664392;
                10'd171  : value <= 32'h3f66894a;
                10'd172  : value <= 32'h3f66cf41;
                10'd173  : value <= 32'h3f671576;
                10'd174  : value <= 32'h3f675be9;
                10'd175  : value <= 32'h3f67a298;
                10'd176  : value <= 32'h3f67e984;
                10'd177  : value <= 32'h3f6830ab;
                10'd178  : value <= 32'h3f68780d;
                10'd179  : value <= 32'h3f68bfaa;
                10'd180  : value <= 32'h3f69077f;
                10'd181  : value <= 32'h3f694f8e;
                10'd182  : value <= 32'h3f6997d5;
                10'd183  : value <= 32'h3f69e053;
                10'd184  : value <= 32'h3f6a2908;
                10'd185  : value <= 32'h3f6a71f2;
                10'd186  : value <= 32'h3f6abb13;
                10'd187  : value <= 32'h3f6b0467;
                10'd188  : value <= 32'h3f6b4df0;
                10'd189  : value <= 32'h3f6b97ab;
                10'd190  : value <= 32'h3f6be19a;
                10'd191  : value <= 32'h3f6c2bb9;
                10'd192  : value <= 32'h3f6c760a;
                10'd193  : value <= 32'h3f6cc08c;
                10'd194  : value <= 32'h3f6d0b3c;
                10'd195  : value <= 32'h3f6d561c;
                10'd196  : value <= 32'h3f6da12a;
                10'd197  : value <= 32'h3f6dec65;
                10'd198  : value <= 32'h3f6e37cd;
                10'd199  : value <= 32'h3f6e8361;
                10'd200  : value <= 32'h3f6ecf20;
                10'd201  : value <= 32'h3f6f1b0a;
                10'd202  : value <= 32'h3f6f671d;
                10'd203  : value <= 32'h3f6fb359;
                10'd204  : value <= 32'h3f6fffbe;
                10'd205  : value <= 32'h3f704c4a;
                10'd206  : value <= 32'h3f7098fd;
                10'd207  : value <= 32'h3f70e5d6;
                10'd208  : value <= 32'h3f7132d5;
                10'd209  : value <= 32'h3f717ff8;
                10'd210  : value <= 32'h3f71cd3f;
                10'd211  : value <= 32'h3f721aa9;
                10'd212  : value <= 32'h3f726835;
                10'd213  : value <= 32'h3f72b5e3;
                10'd214  : value <= 32'h3f7303b2;
                10'd215  : value <= 32'h3f7351a1;
                10'd216  : value <= 32'h3f739faf;
                10'd217  : value <= 32'h3f73eddc;
                10'd218  : value <= 32'h3f743c27;
                10'd219  : value <= 32'h3f748a8f;
                10'd220  : value <= 32'h3f74d913;
                10'd221  : value <= 32'h3f7527b3;
                10'd222  : value <= 32'h3f75766d;
                10'd223  : value <= 32'h3f75c542;
                10'd224  : value <= 32'h3f761430;
                10'd225  : value <= 32'h3f766336;
                10'd226  : value <= 32'h3f76b254;
                10'd227  : value <= 32'h3f770189;
                10'd228  : value <= 32'h3f7750d5;
                10'd229  : value <= 32'h3f77a036;
                10'd230  : value <= 32'h3f77efab;
                10'd231  : value <= 32'h3f783f35;
                10'd232  : value <= 32'h3f788ed1;
                10'd233  : value <= 32'h3f78de80;
                10'd234  : value <= 32'h3f792e41;
                10'd235  : value <= 32'h3f797e13;
                10'd236  : value <= 32'h3f79cdf4;
                10'd237  : value <= 32'h3f7a1de5;
                10'd238  : value <= 32'h3f7a6de5;
                10'd239  : value <= 32'h3f7abdf2;
                10'd240  : value <= 32'h3f7b0e0c;
                10'd241  : value <= 32'h3f7b5e33;
                10'd242  : value <= 32'h3f7bae65;
                10'd243  : value <= 32'h3f7bfea1;
                10'd244  : value <= 32'h3f7c4ee8;
                10'd245  : value <= 32'h3f7c9f38;
                10'd246  : value <= 32'h3f7cef90;
                10'd247  : value <= 32'h3f7d3fef;
                10'd248  : value <= 32'h3f7d9056;
                10'd249  : value <= 32'h3f7de0c2;
                10'd250  : value <= 32'h3f7e3134;
                10'd251  : value <= 32'h3f7e81aa;
                10'd252  : value <= 32'h3f7ed224;
                10'd253  : value <= 32'h3f7f22a0;
                10'd254  : value <= 32'h3f7f731f;
                10'd255  : value <= 32'h3f7fc39f;
                10'd256  : value <= 32'h3f800a10;
                10'd257  : value <= 32'h3f803250;
                10'd258  : value <= 32'h3f805a90;
                10'd259  : value <= 32'h3f8082cf;
                10'd260  : value <= 32'h3f80ab0d;
                10'd261  : value <= 32'h3f80d349;
                10'd262  : value <= 32'h3f80fb83;
                10'd263  : value <= 32'h3f8123ba;
                10'd264  : value <= 32'h3f814bef;
                10'd265  : value <= 32'h3f817421;
                10'd266  : value <= 32'h3f819c4f;
                10'd267  : value <= 32'h3f81c479;
                10'd268  : value <= 32'h3f81ec9e;
                10'd269  : value <= 32'h3f8214bf;
                10'd270  : value <= 32'h3f823cdb;
                10'd271  : value <= 32'h3f8264f1;
                10'd272  : value <= 32'h3f828d01;
                10'd273  : value <= 32'h3f82b50b;
                10'd274  : value <= 32'h3f82dd0e;
                10'd275  : value <= 32'h3f83050b;
                10'd276  : value <= 32'h3f832cff;
                10'd277  : value <= 32'h3f8354ec;
                10'd278  : value <= 32'h3f837cd1;
                10'd279  : value <= 32'h3f83a4ad;
                10'd280  : value <= 32'h3f83cc80;
                10'd281  : value <= 32'h3f83f449;
                10'd282  : value <= 32'h3f841c09;
                10'd283  : value <= 32'h3f8443bf;
                10'd284  : value <= 32'h3f846b6a;
                10'd285  : value <= 32'h3f84930a;
                10'd286  : value <= 32'h3f84ba9f;
                10'd287  : value <= 32'h3f84e228;
                10'd288  : value <= 32'h3f8509a5;
                10'd289  : value <= 32'h3f853116;
                10'd290  : value <= 32'h3f85587a;
                10'd291  : value <= 32'h3f857fd0;
                10'd292  : value <= 32'h3f85a719;
                10'd293  : value <= 32'h3f85ce54;
                10'd294  : value <= 32'h3f85f581;
                10'd295  : value <= 32'h3f861c9f;
                10'd296  : value <= 32'h3f8643ae;
                10'd297  : value <= 32'h3f866aad;
                10'd298  : value <= 32'h3f86919d;
                10'd299  : value <= 32'h3f86b87c;
                10'd300  : value <= 32'h3f86df4b;
                10'd301  : value <= 32'h3f870608;
                10'd302  : value <= 32'h3f872cb4;
                10'd303  : value <= 32'h3f87534f;
                10'd304  : value <= 32'h3f8779d7;
                10'd305  : value <= 32'h3f87a04d;
                10'd306  : value <= 32'h3f87c6b1;
                10'd307  : value <= 32'h3f87ed00;
                10'd308  : value <= 32'h3f88133d;
                10'd309  : value <= 32'h3f883965;
                10'd310  : value <= 32'h3f885f79;
                10'd311  : value <= 32'h3f888578;
                10'd312  : value <= 32'h3f88ab62;
                10'd313  : value <= 32'h3f88d137;
                10'd314  : value <= 32'h3f88f6f6;
                10'd315  : value <= 32'h3f891c9f;
                10'd316  : value <= 32'h3f894231;
                10'd317  : value <= 32'h3f8967ad;
                10'd318  : value <= 32'h3f898d11;
                10'd319  : value <= 32'h3f89b25e;
                10'd320  : value <= 32'h3f89d792;
                10'd321  : value <= 32'h3f89fcae;
                10'd322  : value <= 32'h3f8a21b2;
                10'd323  : value <= 32'h3f8a469c;
                10'd324  : value <= 32'h3f8a6b6d;
                10'd325  : value <= 32'h3f8a9025;
                10'd326  : value <= 32'h3f8ab4c2;
                10'd327  : value <= 32'h3f8ad945;
                10'd328  : value <= 32'h3f8afdad;
                10'd329  : value <= 32'h3f8b21fa;
                10'd330  : value <= 32'h3f8b462b;
                10'd331  : value <= 32'h3f8b6a40;
                10'd332  : value <= 32'h3f8b8e39;
                10'd333  : value <= 32'h3f8bb216;
                10'd334  : value <= 32'h3f8bd5d6;
                10'd335  : value <= 32'h3f8bf978;
                10'd336  : value <= 32'h3f8c1cfd;
                10'd337  : value <= 32'h3f8c4064;
                10'd338  : value <= 32'h3f8c63ac;
                10'd339  : value <= 32'h3f8c86d6;
                10'd340  : value <= 32'h3f8ca9e1;
                10'd341  : value <= 32'h3f8ccccd;
                10'd342  : value <= 32'h3f8cef99;
                10'd343  : value <= 32'h3f8d1245;
                10'd344  : value <= 32'h3f8d34d1;
                10'd345  : value <= 32'h3f8d573c;
                10'd346  : value <= 32'h3f8d7986;
                10'd347  : value <= 32'h3f8d9baf;
                10'd348  : value <= 32'h3f8dbdb6;
                10'd349  : value <= 32'h3f8ddf9b;
                10'd350  : value <= 32'h3f8e015e;
                10'd351  : value <= 32'h3f8e22fe;
                10'd352  : value <= 32'h3f8e447b;
                10'd353  : value <= 32'h3f8e65d5;
                10'd354  : value <= 32'h3f8e870c;
                10'd355  : value <= 32'h3f8ea81e;
                10'd356  : value <= 32'h3f8ec90d;
                10'd357  : value <= 32'h3f8ee9d6;
                10'd358  : value <= 32'h3f8f0a7b;
                10'd359  : value <= 32'h3f8f2afb;
                10'd360  : value <= 32'h3f8f4b55;
                10'd361  : value <= 32'h3f8f6b89;
                10'd362  : value <= 32'h3f8f8b98;
                10'd363  : value <= 32'h3f8fab7f;
                10'd364  : value <= 32'h3f8fcb41;
                10'd365  : value <= 32'h3f8feadb;
                10'd366  : value <= 32'h3f900a4d;
                10'd367  : value <= 32'h3f902998;
                10'd368  : value <= 32'h3f9048bb;
                10'd369  : value <= 32'h3f9067b6;
                10'd370  : value <= 32'h3f908688;
                10'd371  : value <= 32'h3f90a532;
                10'd372  : value <= 32'h3f90c3b2;
                10'd373  : value <= 32'h3f90e209;
                10'd374  : value <= 32'h3f910036;
                10'd375  : value <= 32'h3f911e39;
                10'd376  : value <= 32'h3f913c12;
                10'd377  : value <= 32'h3f9159c0;
                10'd378  : value <= 32'h3f917743;
                10'd379  : value <= 32'h3f91949b;
                10'd380  : value <= 32'h3f91b1c8;
                10'd381  : value <= 32'h3f91cec8;
                10'd382  : value <= 32'h3f91eb9d;
                10'd383  : value <= 32'h3f920846;
                10'd384  : value <= 32'h3f9224c2;
                10'd385  : value <= 32'h3f924111;
                10'd386  : value <= 32'h3f925d33;
                10'd387  : value <= 32'h3f927927;
                10'd388  : value <= 32'h3f9294ee;
                10'd389  : value <= 32'h3f92b087;
                10'd390  : value <= 32'h3f92cbf2;
                10'd391  : value <= 32'h3f92e72e;
                10'd392  : value <= 32'h3f93023b;
                10'd393  : value <= 32'h3f931d1a;
                10'd394  : value <= 32'h3f9337c9;
                10'd395  : value <= 32'h3f935249;
                10'd396  : value <= 32'h3f936c99;
                10'd397  : value <= 32'h3f9386b9;
                10'd398  : value <= 32'h3f93a0a9;
                10'd399  : value <= 32'h3f93ba68;
                10'd400  : value <= 32'h3f93d3f6;
                10'd401  : value <= 32'h3f93ed54;
                10'd402  : value <= 32'h3f940680;
                10'd403  : value <= 32'h3f941f7a;
                10'd404  : value <= 32'h3f943843;
                10'd405  : value <= 32'h3f9450da;
                10'd406  : value <= 32'h3f94693f;
                10'd407  : value <= 32'h3f948171;
                10'd408  : value <= 32'h3f949970;
                10'd409  : value <= 32'h3f94b13d;
                10'd410  : value <= 32'h3f94c8d6;
                10'd411  : value <= 32'h3f94e03c;
                10'd412  : value <= 32'h3f94f76f;
                10'd413  : value <= 32'h3f950e6d;
                10'd414  : value <= 32'h3f952538;
                10'd415  : value <= 32'h3f953bce;
                10'd416  : value <= 32'h3f955230;
                10'd417  : value <= 32'h3f95685d;
                10'd418  : value <= 32'h3f957e55;
                10'd419  : value <= 32'h3f959418;
                10'd420  : value <= 32'h3f95a9a6;
                10'd421  : value <= 32'h3f95befe;
                10'd422  : value <= 32'h3f95d420;
                10'd423  : value <= 32'h3f95e90c;
                10'd424  : value <= 32'h3f95fdc3;
                10'd425  : value <= 32'h3f961242;
                10'd426  : value <= 32'h3f96268c;
                10'd427  : value <= 32'h3f963a9e;
                10'd428  : value <= 32'h3f964e7a;
                10'd429  : value <= 32'h3f96621e;
                10'd430  : value <= 32'h3f96758b;
                10'd431  : value <= 32'h3f9688c1;
                10'd432  : value <= 32'h3f969bbf;
                10'd433  : value <= 32'h3f96ae85;
                10'd434  : value <= 32'h3f96c112;
                10'd435  : value <= 32'h3f96d368;
                10'd436  : value <= 32'h3f96e585;
                10'd437  : value <= 32'h3f96f76a;
                10'd438  : value <= 32'h3f970916;
                10'd439  : value <= 32'h3f971a88;
                10'd440  : value <= 32'h3f972bc2;
                10'd441  : value <= 32'h3f973cc3;
                10'd442  : value <= 32'h3f974d8a;
                10'd443  : value <= 32'h3f975e17;
                10'd444  : value <= 32'h3f976e6b;
                10'd445  : value <= 32'h3f977e84;
                10'd446  : value <= 32'h3f978e64;
                10'd447  : value <= 32'h3f979e09;
                10'd448  : value <= 32'h3f97ad74;
                10'd449  : value <= 32'h3f97bca5;
                10'd450  : value <= 32'h3f97cb9a;
                10'd451  : value <= 32'h3f97da55;
                10'd452  : value <= 32'h3f97e8d5;
                10'd453  : value <= 32'h3f97f71a;
                10'd454  : value <= 32'h3f980524;
                10'd455  : value <= 32'h3f9812f2;
                10'd456  : value <= 32'h3f982085;
                10'd457  : value <= 32'h3f982ddc;
                10'd458  : value <= 32'h3f983af7;
                10'd459  : value <= 32'h3f9847d7;
                10'd460  : value <= 32'h3f98547a;
                10'd461  : value <= 32'h3f9860e1;
                10'd462  : value <= 32'h3f986d0c;
                10'd463  : value <= 32'h3f9878fb;
                10'd464  : value <= 32'h3f9884ad;
                10'd465  : value <= 32'h3f989022;
                10'd466  : value <= 32'h3f989b5b;
                10'd467  : value <= 32'h3f98a657;
                10'd468  : value <= 32'h3f98b116;
                10'd469  : value <= 32'h3f98bb98;
                10'd470  : value <= 32'h3f98c5dc;
                10'd471  : value <= 32'h3f98cfe4;
                10'd472  : value <= 32'h3f98d9ae;
                10'd473  : value <= 32'h3f98e33b;
                10'd474  : value <= 32'h3f98ec8a;
                10'd475  : value <= 32'h3f98f59b;
                10'd476  : value <= 32'h3f98fe6f;
                10'd477  : value <= 32'h3f990705;
                10'd478  : value <= 32'h3f990f5e;
                10'd479  : value <= 32'h3f991778;
                10'd480  : value <= 32'h3f991f54;
                10'd481  : value <= 32'h3f9926f2;
                10'd482  : value <= 32'h3f992e52;
                10'd483  : value <= 32'h3f993574;
                10'd484  : value <= 32'h3f993c57;
                10'd485  : value <= 32'h3f9942fc;
                10'd486  : value <= 32'h3f994963;
                10'd487  : value <= 32'h3f994f8b;
                10'd488  : value <= 32'h3f995574;
                10'd489  : value <= 32'h3f995b1f;
                10'd490  : value <= 32'h3f99608b;
                10'd491  : value <= 32'h3f9965b9;
                10'd492  : value <= 32'h3f996aa7;
                10'd493  : value <= 32'h3f996f57;
                10'd494  : value <= 32'h3f9973c8;
                10'd495  : value <= 32'h3f9977fa;
                10'd496  : value <= 32'h3f997bed;
                10'd497  : value <= 32'h3f997fa1;
                10'd498  : value <= 32'h3f998316;
                10'd499  : value <= 32'h3f99864c;
                10'd500  : value <= 32'h3f998942;
                10'd501  : value <= 32'h3f998bfa;
                10'd502  : value <= 32'h3f998e72;
                10'd503  : value <= 32'h3f9990ac;
                10'd504  : value <= 32'h3f9992a6;
                10'd505  : value <= 32'h3f999461;
                10'd506  : value <= 32'h3f9995dc;
                10'd507  : value <= 32'h3f999719;
                10'd508  : value <= 32'h3f999816;
                10'd509  : value <= 32'h3f9998d4;
                10'd510  : value <= 32'h3f999952;
                10'd511  : value <= 32'h3f999992;
                10'd512  : value <= 32'h3f999992;
                10'd513  : value <= 32'h3f999952;
                10'd514  : value <= 32'h3f9998d4;
                10'd515  : value <= 32'h3f999816;
                10'd516  : value <= 32'h3f999719;
                10'd517  : value <= 32'h3f9995dc;
                10'd518  : value <= 32'h3f999461;
                10'd519  : value <= 32'h3f9992a6;
                10'd520  : value <= 32'h3f9990ac;
                10'd521  : value <= 32'h3f998e72;
                10'd522  : value <= 32'h3f998bfa;
                10'd523  : value <= 32'h3f998942;
                10'd524  : value <= 32'h3f99864c;
                10'd525  : value <= 32'h3f998316;
                10'd526  : value <= 32'h3f997fa1;
                10'd527  : value <= 32'h3f997bed;
                10'd528  : value <= 32'h3f9977fa;
                10'd529  : value <= 32'h3f9973c8;
                10'd530  : value <= 32'h3f996f57;
                10'd531  : value <= 32'h3f996aa7;
                10'd532  : value <= 32'h3f9965b9;
                10'd533  : value <= 32'h3f99608b;
                10'd534  : value <= 32'h3f995b1f;
                10'd535  : value <= 32'h3f995574;
                10'd536  : value <= 32'h3f994f8b;
                10'd537  : value <= 32'h3f994963;
                10'd538  : value <= 32'h3f9942fc;
                10'd539  : value <= 32'h3f993c57;
                10'd540  : value <= 32'h3f993574;
                10'd541  : value <= 32'h3f992e52;
                10'd542  : value <= 32'h3f9926f2;
                10'd543  : value <= 32'h3f991f54;
                10'd544  : value <= 32'h3f991778;
                10'd545  : value <= 32'h3f990f5e;
                10'd546  : value <= 32'h3f990705;
                10'd547  : value <= 32'h3f98fe6f;
                10'd548  : value <= 32'h3f98f59b;
                10'd549  : value <= 32'h3f98ec8a;
                10'd550  : value <= 32'h3f98e33b;
                10'd551  : value <= 32'h3f98d9ae;
                10'd552  : value <= 32'h3f98cfe4;
                10'd553  : value <= 32'h3f98c5dc;
                10'd554  : value <= 32'h3f98bb98;
                10'd555  : value <= 32'h3f98b116;
                10'd556  : value <= 32'h3f98a657;
                10'd557  : value <= 32'h3f989b5b;
                10'd558  : value <= 32'h3f989022;
                10'd559  : value <= 32'h3f9884ad;
                10'd560  : value <= 32'h3f9878fb;
                10'd561  : value <= 32'h3f986d0c;
                10'd562  : value <= 32'h3f9860e1;
                10'd563  : value <= 32'h3f98547a;
                10'd564  : value <= 32'h3f9847d7;
                10'd565  : value <= 32'h3f983af7;
                10'd566  : value <= 32'h3f982ddc;
                10'd567  : value <= 32'h3f982085;
                10'd568  : value <= 32'h3f9812f2;
                10'd569  : value <= 32'h3f980524;
                10'd570  : value <= 32'h3f97f71a;
                10'd571  : value <= 32'h3f97e8d5;
                10'd572  : value <= 32'h3f97da55;
                10'd573  : value <= 32'h3f97cb9a;
                10'd574  : value <= 32'h3f97bca5;
                10'd575  : value <= 32'h3f97ad74;
                10'd576  : value <= 32'h3f979e09;
                10'd577  : value <= 32'h3f978e64;
                10'd578  : value <= 32'h3f977e84;
                10'd579  : value <= 32'h3f976e6b;
                10'd580  : value <= 32'h3f975e17;
                10'd581  : value <= 32'h3f974d8a;
                10'd582  : value <= 32'h3f973cc3;
                10'd583  : value <= 32'h3f972bc2;
                10'd584  : value <= 32'h3f971a88;
                10'd585  : value <= 32'h3f970916;
                10'd586  : value <= 32'h3f96f76a;
                10'd587  : value <= 32'h3f96e585;
                10'd588  : value <= 32'h3f96d368;
                10'd589  : value <= 32'h3f96c112;
                10'd590  : value <= 32'h3f96ae85;
                10'd591  : value <= 32'h3f969bbf;
                10'd592  : value <= 32'h3f9688c1;
                10'd593  : value <= 32'h3f96758b;
                10'd594  : value <= 32'h3f96621e;
                10'd595  : value <= 32'h3f964e7a;
                10'd596  : value <= 32'h3f963a9e;
                10'd597  : value <= 32'h3f96268c;
                10'd598  : value <= 32'h3f961242;
                10'd599  : value <= 32'h3f95fdc3;
                10'd600  : value <= 32'h3f95e90c;
                10'd601  : value <= 32'h3f95d420;
                10'd602  : value <= 32'h3f95befe;
                10'd603  : value <= 32'h3f95a9a6;
                10'd604  : value <= 32'h3f959418;
                10'd605  : value <= 32'h3f957e55;
                10'd606  : value <= 32'h3f95685d;
                10'd607  : value <= 32'h3f955230;
                10'd608  : value <= 32'h3f953bce;
                10'd609  : value <= 32'h3f952538;
                10'd610  : value <= 32'h3f950e6d;
                10'd611  : value <= 32'h3f94f76f;
                10'd612  : value <= 32'h3f94e03c;
                10'd613  : value <= 32'h3f94c8d6;
                10'd614  : value <= 32'h3f94b13d;
                10'd615  : value <= 32'h3f949970;
                10'd616  : value <= 32'h3f948171;
                10'd617  : value <= 32'h3f94693f;
                10'd618  : value <= 32'h3f9450da;
                10'd619  : value <= 32'h3f943843;
                10'd620  : value <= 32'h3f941f7a;
                10'd621  : value <= 32'h3f940680;
                10'd622  : value <= 32'h3f93ed54;
                10'd623  : value <= 32'h3f93d3f6;
                10'd624  : value <= 32'h3f93ba68;
                10'd625  : value <= 32'h3f93a0a9;
                10'd626  : value <= 32'h3f9386b9;
                10'd627  : value <= 32'h3f936c99;
                10'd628  : value <= 32'h3f935249;
                10'd629  : value <= 32'h3f9337c9;
                10'd630  : value <= 32'h3f931d1a;
                10'd631  : value <= 32'h3f93023b;
                10'd632  : value <= 32'h3f92e72e;
                10'd633  : value <= 32'h3f92cbf2;
                10'd634  : value <= 32'h3f92b087;
                10'd635  : value <= 32'h3f9294ee;
                10'd636  : value <= 32'h3f927927;
                10'd637  : value <= 32'h3f925d33;
                10'd638  : value <= 32'h3f924111;
                10'd639  : value <= 32'h3f9224c2;
                10'd640  : value <= 32'h3f920846;
                10'd641  : value <= 32'h3f91eb9d;
                10'd642  : value <= 32'h3f91cec8;
                10'd643  : value <= 32'h3f91b1c8;
                10'd644  : value <= 32'h3f91949b;
                10'd645  : value <= 32'h3f917743;
                10'd646  : value <= 32'h3f9159c0;
                10'd647  : value <= 32'h3f913c12;
                10'd648  : value <= 32'h3f911e39;
                10'd649  : value <= 32'h3f910036;
                10'd650  : value <= 32'h3f90e209;
                10'd651  : value <= 32'h3f90c3b2;
                10'd652  : value <= 32'h3f90a532;
                10'd653  : value <= 32'h3f908688;
                10'd654  : value <= 32'h3f9067b6;
                10'd655  : value <= 32'h3f9048bb;
                10'd656  : value <= 32'h3f902998;
                10'd657  : value <= 32'h3f900a4d;
                10'd658  : value <= 32'h3f8feadb;
                10'd659  : value <= 32'h3f8fcb41;
                10'd660  : value <= 32'h3f8fab7f;
                10'd661  : value <= 32'h3f8f8b98;
                10'd662  : value <= 32'h3f8f6b89;
                10'd663  : value <= 32'h3f8f4b55;
                10'd664  : value <= 32'h3f8f2afb;
                10'd665  : value <= 32'h3f8f0a7b;
                10'd666  : value <= 32'h3f8ee9d6;
                10'd667  : value <= 32'h3f8ec90d;
                10'd668  : value <= 32'h3f8ea81e;
                10'd669  : value <= 32'h3f8e870c;
                10'd670  : value <= 32'h3f8e65d5;
                10'd671  : value <= 32'h3f8e447b;
                10'd672  : value <= 32'h3f8e22fe;
                10'd673  : value <= 32'h3f8e015e;
                10'd674  : value <= 32'h3f8ddf9b;
                10'd675  : value <= 32'h3f8dbdb6;
                10'd676  : value <= 32'h3f8d9baf;
                10'd677  : value <= 32'h3f8d7986;
                10'd678  : value <= 32'h3f8d573c;
                10'd679  : value <= 32'h3f8d34d1;
                10'd680  : value <= 32'h3f8d1245;
                10'd681  : value <= 32'h3f8cef99;
                10'd682  : value <= 32'h3f8ccccd;
                10'd683  : value <= 32'h3f8ca9e1;
                10'd684  : value <= 32'h3f8c86d6;
                10'd685  : value <= 32'h3f8c63ac;
                10'd686  : value <= 32'h3f8c4064;
                10'd687  : value <= 32'h3f8c1cfd;
                10'd688  : value <= 32'h3f8bf978;
                10'd689  : value <= 32'h3f8bd5d6;
                10'd690  : value <= 32'h3f8bb216;
                10'd691  : value <= 32'h3f8b8e39;
                10'd692  : value <= 32'h3f8b6a40;
                10'd693  : value <= 32'h3f8b462b;
                10'd694  : value <= 32'h3f8b21fa;
                10'd695  : value <= 32'h3f8afdad;
                10'd696  : value <= 32'h3f8ad945;
                10'd697  : value <= 32'h3f8ab4c2;
                10'd698  : value <= 32'h3f8a9025;
                10'd699  : value <= 32'h3f8a6b6d;
                10'd700  : value <= 32'h3f8a469c;
                10'd701  : value <= 32'h3f8a21b2;
                10'd702  : value <= 32'h3f89fcae;
                10'd703  : value <= 32'h3f89d792;
                10'd704  : value <= 32'h3f89b25e;
                10'd705  : value <= 32'h3f898d11;
                10'd706  : value <= 32'h3f8967ad;
                10'd707  : value <= 32'h3f894231;
                10'd708  : value <= 32'h3f891c9f;
                10'd709  : value <= 32'h3f88f6f6;
                10'd710  : value <= 32'h3f88d137;
                10'd711  : value <= 32'h3f88ab62;
                10'd712  : value <= 32'h3f888578;
                10'd713  : value <= 32'h3f885f79;
                10'd714  : value <= 32'h3f883965;
                10'd715  : value <= 32'h3f88133d;
                10'd716  : value <= 32'h3f87ed00;
                10'd717  : value <= 32'h3f87c6b1;
                10'd718  : value <= 32'h3f87a04d;
                10'd719  : value <= 32'h3f8779d7;
                10'd720  : value <= 32'h3f87534f;
                10'd721  : value <= 32'h3f872cb4;
                10'd722  : value <= 32'h3f870608;
                10'd723  : value <= 32'h3f86df4b;
                10'd724  : value <= 32'h3f86b87c;
                10'd725  : value <= 32'h3f86919d;
                10'd726  : value <= 32'h3f866aad;
                10'd727  : value <= 32'h3f8643ae;
                10'd728  : value <= 32'h3f861c9f;
                10'd729  : value <= 32'h3f85f581;
                10'd730  : value <= 32'h3f85ce54;
                10'd731  : value <= 32'h3f85a719;
                10'd732  : value <= 32'h3f857fd0;
                10'd733  : value <= 32'h3f85587a;
                10'd734  : value <= 32'h3f853116;
                10'd735  : value <= 32'h3f8509a5;
                10'd736  : value <= 32'h3f84e228;
                10'd737  : value <= 32'h3f84ba9f;
                10'd738  : value <= 32'h3f84930a;
                10'd739  : value <= 32'h3f846b6a;
                10'd740  : value <= 32'h3f8443bf;
                10'd741  : value <= 32'h3f841c09;
                10'd742  : value <= 32'h3f83f449;
                10'd743  : value <= 32'h3f83cc80;
                10'd744  : value <= 32'h3f83a4ad;
                10'd745  : value <= 32'h3f837cd1;
                10'd746  : value <= 32'h3f8354ec;
                10'd747  : value <= 32'h3f832cff;
                10'd748  : value <= 32'h3f83050b;
                10'd749  : value <= 32'h3f82dd0e;
                10'd750  : value <= 32'h3f82b50b;
                10'd751  : value <= 32'h3f828d01;
                10'd752  : value <= 32'h3f8264f1;
                10'd753  : value <= 32'h3f823cdb;
                10'd754  : value <= 32'h3f8214bf;
                10'd755  : value <= 32'h3f81ec9e;
                10'd756  : value <= 32'h3f81c479;
                10'd757  : value <= 32'h3f819c4f;
                10'd758  : value <= 32'h3f817421;
                10'd759  : value <= 32'h3f814bef;
                10'd760  : value <= 32'h3f8123ba;
                10'd761  : value <= 32'h3f80fb83;
                10'd762  : value <= 32'h3f80d349;
                10'd763  : value <= 32'h3f80ab0d;
                10'd764  : value <= 32'h3f8082cf;
                10'd765  : value <= 32'h3f805a90;
                10'd766  : value <= 32'h3f803250;
                10'd767  : value <= 32'h3f800a10;
                10'd768  : value <= 32'h3f7fc39f;
                10'd769  : value <= 32'h3f7f731f;
                10'd770  : value <= 32'h3f7f22a0;
                10'd771  : value <= 32'h3f7ed224;
                10'd772  : value <= 32'h3f7e81aa;
                10'd773  : value <= 32'h3f7e3134;
                10'd774  : value <= 32'h3f7de0c2;
                10'd775  : value <= 32'h3f7d9056;
                10'd776  : value <= 32'h3f7d3fef;
                10'd777  : value <= 32'h3f7cef90;
                10'd778  : value <= 32'h3f7c9f38;
                10'd779  : value <= 32'h3f7c4ee8;
                10'd780  : value <= 32'h3f7bfea1;
                10'd781  : value <= 32'h3f7bae65;
                10'd782  : value <= 32'h3f7b5e33;
                10'd783  : value <= 32'h3f7b0e0c;
                10'd784  : value <= 32'h3f7abdf2;
                10'd785  : value <= 32'h3f7a6de5;
                10'd786  : value <= 32'h3f7a1de5;
                10'd787  : value <= 32'h3f79cdf4;
                10'd788  : value <= 32'h3f797e13;
                10'd789  : value <= 32'h3f792e41;
                10'd790  : value <= 32'h3f78de80;
                10'd791  : value <= 32'h3f788ed1;
                10'd792  : value <= 32'h3f783f35;
                10'd793  : value <= 32'h3f77efab;
                10'd794  : value <= 32'h3f77a036;
                10'd795  : value <= 32'h3f7750d5;
                10'd796  : value <= 32'h3f770189;
                10'd797  : value <= 32'h3f76b254;
                10'd798  : value <= 32'h3f766336;
                10'd799  : value <= 32'h3f761430;
                10'd800  : value <= 32'h3f75c542;
                10'd801  : value <= 32'h3f75766d;
                10'd802  : value <= 32'h3f7527b3;
                10'd803  : value <= 32'h3f74d913;
                10'd804  : value <= 32'h3f748a8f;
                10'd805  : value <= 32'h3f743c27;
                10'd806  : value <= 32'h3f73eddc;
                10'd807  : value <= 32'h3f739faf;
                10'd808  : value <= 32'h3f7351a1;
                10'd809  : value <= 32'h3f7303b2;
                10'd810  : value <= 32'h3f72b5e3;
                10'd811  : value <= 32'h3f726835;
                10'd812  : value <= 32'h3f721aa9;
                10'd813  : value <= 32'h3f71cd3f;
                10'd814  : value <= 32'h3f717ff8;
                10'd815  : value <= 32'h3f7132d5;
                10'd816  : value <= 32'h3f70e5d6;
                10'd817  : value <= 32'h3f7098fd;
                10'd818  : value <= 32'h3f704c4a;
                10'd819  : value <= 32'h3f6fffbe;
                10'd820  : value <= 32'h3f6fb359;
                10'd821  : value <= 32'h3f6f671d;
                10'd822  : value <= 32'h3f6f1b0a;
                10'd823  : value <= 32'h3f6ecf20;
                10'd824  : value <= 32'h3f6e8361;
                10'd825  : value <= 32'h3f6e37cd;
                10'd826  : value <= 32'h3f6dec65;
                10'd827  : value <= 32'h3f6da12a;
                10'd828  : value <= 32'h3f6d561c;
                10'd829  : value <= 32'h3f6d0b3c;
                10'd830  : value <= 32'h3f6cc08c;
                10'd831  : value <= 32'h3f6c760a;
                10'd832  : value <= 32'h3f6c2bb9;
                10'd833  : value <= 32'h3f6be19a;
                10'd834  : value <= 32'h3f6b97ab;
                10'd835  : value <= 32'h3f6b4df0;
                10'd836  : value <= 32'h3f6b0467;
                10'd837  : value <= 32'h3f6abb13;
                10'd838  : value <= 32'h3f6a71f2;
                10'd839  : value <= 32'h3f6a2908;
                10'd840  : value <= 32'h3f69e053;
                10'd841  : value <= 32'h3f6997d5;
                10'd842  : value <= 32'h3f694f8e;
                10'd843  : value <= 32'h3f69077f;
                10'd844  : value <= 32'h3f68bfaa;
                10'd845  : value <= 32'h3f68780d;
                10'd846  : value <= 32'h3f6830ab;
                10'd847  : value <= 32'h3f67e984;
                10'd848  : value <= 32'h3f67a298;
                10'd849  : value <= 32'h3f675be9;
                10'd850  : value <= 32'h3f671576;
                10'd851  : value <= 32'h3f66cf41;
                10'd852  : value <= 32'h3f66894a;
                10'd853  : value <= 32'h3f664392;
                10'd854  : value <= 32'h3f65fe1a;
                10'd855  : value <= 32'h3f65b8e2;
                10'd856  : value <= 32'h3f6573ec;
                10'd857  : value <= 32'h3f652f36;
                10'd858  : value <= 32'h3f64eac3;
                10'd859  : value <= 32'h3f64a693;
                10'd860  : value <= 32'h3f6462a7;
                10'd861  : value <= 32'h3f641eff;
                10'd862  : value <= 32'h3f63db9c;
                10'd863  : value <= 32'h3f63987e;
                10'd864  : value <= 32'h3f6355a7;
                10'd865  : value <= 32'h3f631316;
                10'd866  : value <= 32'h3f62d0cd;
                10'd867  : value <= 32'h3f628ecc;
                10'd868  : value <= 32'h3f624d14;
                10'd869  : value <= 32'h3f620ba5;
                10'd870  : value <= 32'h3f61ca81;
                10'd871  : value <= 32'h3f6189a7;
                10'd872  : value <= 32'h3f614918;
                10'd873  : value <= 32'h3f6108d5;
                10'd874  : value <= 32'h3f60c8df;
                10'd875  : value <= 32'h3f608936;
                10'd876  : value <= 32'h3f6049db;
                10'd877  : value <= 32'h3f600ace;
                10'd878  : value <= 32'h3f5fcc11;
                10'd879  : value <= 32'h3f5f8da2;
                10'd880  : value <= 32'h3f5f4f84;
                10'd881  : value <= 32'h3f5f11b7;
                10'd882  : value <= 32'h3f5ed43c;
                10'd883  : value <= 32'h3f5e9712;
                10'd884  : value <= 32'h3f5e5a3b;
                10'd885  : value <= 32'h3f5e1db7;
                10'd886  : value <= 32'h3f5de187;
                10'd887  : value <= 32'h3f5da5ab;
                10'd888  : value <= 32'h3f5d6a24;
                10'd889  : value <= 32'h3f5d2ef3;
                10'd890  : value <= 32'h3f5cf417;
                10'd891  : value <= 32'h3f5cb993;
                10'd892  : value <= 32'h3f5c7f65;
                10'd893  : value <= 32'h3f5c458f;
                10'd894  : value <= 32'h3f5c0c12;
                10'd895  : value <= 32'h3f5bd2ee;
                10'd896  : value <= 32'h3f5b9a23;
                10'd897  : value <= 32'h3f5b61b2;
                10'd898  : value <= 32'h3f5b299b;
                10'd899  : value <= 32'h3f5af1e0;
                10'd900  : value <= 32'h3f5aba80;
                10'd901  : value <= 32'h3f5a837c;
                10'd902  : value <= 32'h3f5a4cd5;
                10'd903  : value <= 32'h3f5a168b;
                10'd904  : value <= 32'h3f59e09f;
                10'd905  : value <= 32'h3f59ab11;
                10'd906  : value <= 32'h3f5975e2;
                10'd907  : value <= 32'h3f594112;
                10'd908  : value <= 32'h3f590ca2;
                10'd909  : value <= 32'h3f58d892;
                10'd910  : value <= 32'h3f58a4e4;
                10'd911  : value <= 32'h3f587196;
                10'd912  : value <= 32'h3f583eaa;
                10'd913  : value <= 32'h3f580c20;
                10'd914  : value <= 32'h3f57d9fa;
                10'd915  : value <= 32'h3f57a836;
                10'd916  : value <= 32'h3f5776d6;
                10'd917  : value <= 32'h3f5745db;
                10'd918  : value <= 32'h3f571544;
                10'd919  : value <= 32'h3f56e512;
                10'd920  : value <= 32'h3f56b546;
                10'd921  : value <= 32'h3f5685e0;
                10'd922  : value <= 32'h3f5656e0;
                10'd923  : value <= 32'h3f562848;
                10'd924  : value <= 32'h3f55fa17;
                10'd925  : value <= 32'h3f55cc4e;
                10'd926  : value <= 32'h3f559eed;
                10'd927  : value <= 32'h3f5571f5;
                10'd928  : value <= 32'h3f554566;
                10'd929  : value <= 32'h3f551941;
                10'd930  : value <= 32'h3f54ed86;
                10'd931  : value <= 32'h3f54c235;
                10'd932  : value <= 32'h3f54974f;
                10'd933  : value <= 32'h3f546cd5;
                10'd934  : value <= 32'h3f5442c6;
                10'd935  : value <= 32'h3f541923;
                10'd936  : value <= 32'h3f53efed;
                10'd937  : value <= 32'h3f53c724;
                10'd938  : value <= 32'h3f539ec8;
                10'd939  : value <= 32'h3f5376da;
                10'd940  : value <= 32'h3f534f5a;
                10'd941  : value <= 32'h3f532849;
                10'd942  : value <= 32'h3f5301a6;
                10'd943  : value <= 32'h3f52db73;
                10'd944  : value <= 32'h3f52b5af;
                10'd945  : value <= 32'h3f52905b;
                10'd946  : value <= 32'h3f526b77;
                10'd947  : value <= 32'h3f524705;
                10'd948  : value <= 32'h3f522303;
                10'd949  : value <= 32'h3f51ff72;
                10'd950  : value <= 32'h3f51dc54;
                10'd951  : value <= 32'h3f51b9a7;
                10'd952  : value <= 32'h3f51976d;
                10'd953  : value <= 32'h3f5175a5;
                10'd954  : value <= 32'h3f515451;
                10'd955  : value <= 32'h3f513370;
                10'd956  : value <= 32'h3f511303;
                10'd957  : value <= 32'h3f50f309;
                10'd958  : value <= 32'h3f50d384;
                10'd959  : value <= 32'h3f50b474;
                10'd960  : value <= 32'h3f5095d8;
                10'd961  : value <= 32'h3f5077b2;
                10'd962  : value <= 32'h3f505a01;
                10'd963  : value <= 32'h3f503cc6;
                10'd964  : value <= 32'h3f502002;
                10'd965  : value <= 32'h3f5003b3;
                10'd966  : value <= 32'h3f4fe7db;
                10'd967  : value <= 32'h3f4fcc7a;
                10'd968  : value <= 32'h3f4fb190;
                10'd969  : value <= 32'h3f4f971e;
                10'd970  : value <= 32'h3f4f7d23;
                10'd971  : value <= 32'h3f4f63a1;
                10'd972  : value <= 32'h3f4f4a96;
                10'd973  : value <= 32'h3f4f3204;
                10'd974  : value <= 32'h3f4f19ea;
                10'd975  : value <= 32'h3f4f024a;
                10'd976  : value <= 32'h3f4eeb22;
                10'd977  : value <= 32'h3f4ed474;
                10'd978  : value <= 32'h3f4ebe3f;
                10'd979  : value <= 32'h3f4ea884;
                10'd980  : value <= 32'h3f4e9344;
                10'd981  : value <= 32'h3f4e7e7d;
                10'd982  : value <= 32'h3f4e6a31;
                10'd983  : value <= 32'h3f4e565f;
                10'd984  : value <= 32'h3f4e4308;
                10'd985  : value <= 32'h3f4e302c;
                10'd986  : value <= 32'h3f4e1dcb;
                10'd987  : value <= 32'h3f4e0be6;
                10'd988  : value <= 32'h3f4dfa7c;
                10'd989  : value <= 32'h3f4de98d;
                10'd990  : value <= 32'h3f4dd91b;
                10'd991  : value <= 32'h3f4dc924;
                10'd992  : value <= 32'h3f4db9aa;
                10'd993  : value <= 32'h3f4daaac;
                10'd994  : value <= 32'h3f4d9c2a;
                10'd995  : value <= 32'h3f4d8e25;
                10'd996  : value <= 32'h3f4d809d;
                10'd997  : value <= 32'h3f4d7391;
                10'd998  : value <= 32'h3f4d6703;
                10'd999  : value <= 32'h3f4d5af1;
                10'd1000  : value <= 32'h3f4d4f5d;
                10'd1001  : value <= 32'h3f4d4446;
                10'd1002  : value <= 32'h3f4d39ad;
                10'd1003  : value <= 32'h3f4d2f91;
                10'd1004  : value <= 32'h3f4d25f2;
                10'd1005  : value <= 32'h3f4d1cd2;
                10'd1006  : value <= 32'h3f4d142f;
                10'd1007  : value <= 32'h3f4d0c0a;
                10'd1008  : value <= 32'h3f4d0463;
                10'd1009  : value <= 32'h3f4cfd3a;
                10'd1010  : value <= 32'h3f4cf68f;
                10'd1011  : value <= 32'h3f4cf062;
                10'd1012  : value <= 32'h3f4ceab4;
                10'd1013  : value <= 32'h3f4ce584;
                10'd1014  : value <= 32'h3f4ce0d2;
                10'd1015  : value <= 32'h3f4cdc9e;
                10'd1016  : value <= 32'h3f4cd8e9;
                10'd1017  : value <= 32'h3f4cd5b3;
                10'd1018  : value <= 32'h3f4cd2fb;
                10'd1019  : value <= 32'h3f4cd0c1;
                10'd1020  : value <= 32'h3f4ccf06;
                10'd1021  : value <= 32'h3f4ccdca;
                10'd1022  : value <= 32'h3f4ccd0c;
                10'd1023  : value <= 32'h3f4ccccd;
                default   : value <= 32'h3f4ccccd;
            endcase
        end // if not reset
    end
endmodule
