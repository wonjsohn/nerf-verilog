`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:04:56 07/18/2011 
// Design Name: 
// Module Name:    spindle_neuron 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module spindle_neuron(	input [31:0] pps,
								input clk,
                        input reset,
								output reg spike
    );

	reg [10:0] isi_count; //Inter spike interval count
	reg [10:0] spike_count;	//spike count over 1 second
	reg [1023:0] spike_history;
    wire [31:0] floored_pps;
	wire [10:0] int_pps;
	wire [10:0] isi;			//inter spike interval based on pps firing rate
	wire [10:0] isi_final;	//inter spike interval taking into account fractional isi
	
	wire generate_spike; //command to spike on this clock cycle
	
    
    floor floor1(.in(pps), .out(floored_pps));
    assign int_pps = floored_pps[10:0];
	 
	pps_to_isi pi_convertor( .pps(int_pps), .isi(isi) );
	
	assign isi_final = (spike_count > int_pps) ? (isi+1) : (isi); //if over-firing, delay spike 1 cycle
	
	assign generate_spike = (isi_count >= isi_final) ? 1'b1 : 1'b0;
	
	always @ (posedge clk)
	begin
		// this section if generate_spike == 0
		isi_count <= isi_count+1;
		spike <= generate_spike;
		spike_history <= {spike_history[1022:0], generate_spike};
		spike_count <= spike_count - spike_history[1023] + generate_spike;
		
		if (reset)
		begin
			//this section on reset
			isi_count <= 1;
			spike_history <= 1023'd0;
			spike <= 0;
			spike_count <= 0;
		end
		else if (generate_spike)
		begin
			//this section if generate_spike == 1
			isi_count <= 1;
			spike_history <= {spike_history[1022:0], generate_spike};
			spike <= generate_spike;
			spike_count <= spike_count - spike_history[1023] + generate_spike;
		end
	end
	
endmodule

module pps_to_isi( 	input [10:0] pps,
							output reg [10:0] isi );
							
//Convert firing rate (pulses per second) to inter-spike interval
//reciprocal function too expensive, use Look-up table

    always @ (pps)
    begin
    case (pps)
                11'd0  : isi = 11'h400;
                11'd1  : isi = 11'h200;
                11'd2  : isi = 11'h155;
                11'd3  : isi = 11'h100;
                11'd4  : isi = 11'hcc;
                11'd5  : isi = 11'haa;
                11'd6  : isi = 11'h92;
                11'd7  : isi = 11'h80;
                11'd8  : isi = 11'h71;
                11'd9  : isi = 11'h66;
                11'd10  : isi = 11'h5d;
                11'd11  : isi = 11'h55;
                11'd12  : isi = 11'h4e;
                11'd13  : isi = 11'h49;
                11'd14  : isi = 11'h44;
                11'd15  : isi = 11'h40;
                11'd16  : isi = 11'h3c;
                11'd17  : isi = 11'h38;
                11'd18  : isi = 11'h35;
                11'd19  : isi = 11'h33;
                11'd20  : isi = 11'h30;
                11'd21  : isi = 11'h2e;
                11'd22  : isi = 11'h2c;
                11'd23  : isi = 11'h2a;
                11'd24  : isi = 11'h28;
                11'd25  : isi = 11'h27;
                11'd26  : isi = 11'h25;
                11'd27  : isi = 11'h24;
                11'd28  : isi = 11'h23;
                11'd29  : isi = 11'h22;
                11'd30  : isi = 11'h21;
                11'd31  : isi = 11'h20;
                11'd32  : isi = 11'h1f;
                11'd33  : isi = 11'h1e;
                11'd34  : isi = 11'h1d;
                11'd35  : isi = 11'h1c;
                11'd36  : isi = 11'h1b;
                11'd37  : isi = 11'h1a;
                11'd38  : isi = 11'h1a;
                11'd39  : isi = 11'h19;
                11'd40  : isi = 11'h18;
                11'd41  : isi = 11'h18;
                11'd42  : isi = 11'h17;
                11'd43  : isi = 11'h17;
                11'd44  : isi = 11'h16;
                11'd45  : isi = 11'h16;
                11'd46  : isi = 11'h15;
                11'd47  : isi = 11'h15;
                11'd48  : isi = 11'h14;
                11'd49  : isi = 11'h14;
                11'd50  : isi = 11'h14;
                11'd51  : isi = 11'h13;
                11'd52  : isi = 11'h13;
                11'd53  : isi = 11'h12;
                11'd54  : isi = 11'h12;
                11'd55  : isi = 11'h12;
                11'd56  : isi = 11'h11;
                11'd57  : isi = 11'h11;
                11'd58  : isi = 11'h11;
                11'd59  : isi = 11'h11;
                11'd60  : isi = 11'h10;
                11'd61  : isi = 11'h10;
                11'd62  : isi = 11'h10;
                11'd63  : isi = 11'h10;
                11'd64  : isi = 11'hf;
                11'd65  : isi = 11'hf;
                11'd66  : isi = 11'hf;
                11'd67  : isi = 11'hf;
                11'd68  : isi = 11'he;
                11'd69  : isi = 11'he;
                11'd70  : isi = 11'he;
                11'd71  : isi = 11'he;
                11'd72  : isi = 11'he;
                11'd73  : isi = 11'hd;
                11'd74  : isi = 11'hd;
                11'd75  : isi = 11'hd;
                11'd76  : isi = 11'hd;
                11'd77  : isi = 11'hd;
                11'd78  : isi = 11'hc;
                11'd79  : isi = 11'hc;
                11'd80  : isi = 11'hc;
                11'd81  : isi = 11'hc;
                11'd82  : isi = 11'hc;
                11'd83  : isi = 11'hc;
                11'd84  : isi = 11'hc;
                11'd85  : isi = 11'hb;
                11'd86  : isi = 11'hb;
                11'd87  : isi = 11'hb;
                11'd88  : isi = 11'hb;
                11'd89  : isi = 11'hb;
                11'd90  : isi = 11'hb;
                11'd91  : isi = 11'hb;
                11'd92  : isi = 11'hb;
                11'd93  : isi = 11'ha;
                11'd94  : isi = 11'ha;
                11'd95  : isi = 11'ha;
                11'd96  : isi = 11'ha;
                11'd97  : isi = 11'ha;
                11'd98  : isi = 11'ha;
                11'd99  : isi = 11'ha;
                11'd100  : isi = 11'ha;
                11'd101  : isi = 11'ha;
                11'd102  : isi = 11'h9;
                11'd103  : isi = 11'h9;
                11'd104  : isi = 11'h9;
                11'd105  : isi = 11'h9;
                11'd106  : isi = 11'h9;
                11'd107  : isi = 11'h9;
                11'd108  : isi = 11'h9;
                11'd109  : isi = 11'h9;
                11'd110  : isi = 11'h9;
                11'd111  : isi = 11'h9;
                11'd112  : isi = 11'h9;
                11'd113  : isi = 11'h8;
                11'd114  : isi = 11'h8;
                11'd115  : isi = 11'h8;
                11'd116  : isi = 11'h8;
                11'd117  : isi = 11'h8;
                11'd118  : isi = 11'h8;
                11'd119  : isi = 11'h8;
                11'd120  : isi = 11'h8;
                11'd121  : isi = 11'h8;
                11'd122  : isi = 11'h8;
                11'd123  : isi = 11'h8;
                11'd124  : isi = 11'h8;
                11'd125  : isi = 11'h8;
                11'd126  : isi = 11'h8;
                11'd127  : isi = 11'h8;
                11'd128  : isi = 11'h7;
                11'd129  : isi = 11'h7;
                11'd130  : isi = 11'h7;
                11'd131  : isi = 11'h7;
                11'd132  : isi = 11'h7;
                11'd133  : isi = 11'h7;
                11'd134  : isi = 11'h7;
                11'd135  : isi = 11'h7;
                11'd136  : isi = 11'h7;
                11'd137  : isi = 11'h7;
                11'd138  : isi = 11'h7;
                11'd139  : isi = 11'h7;
                11'd140  : isi = 11'h7;
                11'd141  : isi = 11'h7;
                11'd142  : isi = 11'h7;
                11'd143  : isi = 11'h7;
                11'd144  : isi = 11'h7;
                11'd145  : isi = 11'h7;
                11'd146  : isi = 11'h6;
                11'd147  : isi = 11'h6;
                11'd148  : isi = 11'h6;
                11'd149  : isi = 11'h6;
                11'd150  : isi = 11'h6;
                11'd151  : isi = 11'h6;
                11'd152  : isi = 11'h6;
                11'd153  : isi = 11'h6;
                11'd154  : isi = 11'h6;
                11'd155  : isi = 11'h6;
                11'd156  : isi = 11'h6;
                11'd157  : isi = 11'h6;
                11'd158  : isi = 11'h6;
                11'd159  : isi = 11'h6;
                11'd160  : isi = 11'h6;
                11'd161  : isi = 11'h6;
                11'd162  : isi = 11'h6;
                11'd163  : isi = 11'h6;
                11'd164  : isi = 11'h6;
                11'd165  : isi = 11'h6;
                11'd166  : isi = 11'h6;
                11'd167  : isi = 11'h6;
                11'd168  : isi = 11'h6;
                11'd169  : isi = 11'h6;
                11'd170  : isi = 11'h5;
                11'd171  : isi = 11'h5;
                11'd172  : isi = 11'h5;
                11'd173  : isi = 11'h5;
                11'd174  : isi = 11'h5;
                11'd175  : isi = 11'h5;
                11'd176  : isi = 11'h5;
                11'd177  : isi = 11'h5;
                11'd178  : isi = 11'h5;
                11'd179  : isi = 11'h5;
                11'd180  : isi = 11'h5;
                11'd181  : isi = 11'h5;
                11'd182  : isi = 11'h5;
                11'd183  : isi = 11'h5;
                11'd184  : isi = 11'h5;
                11'd185  : isi = 11'h5;
                11'd186  : isi = 11'h5;
                11'd187  : isi = 11'h5;
                11'd188  : isi = 11'h5;
                11'd189  : isi = 11'h5;
                11'd190  : isi = 11'h5;
                11'd191  : isi = 11'h5;
                11'd192  : isi = 11'h5;
                11'd193  : isi = 11'h5;
                11'd194  : isi = 11'h5;
                11'd195  : isi = 11'h5;
                11'd196  : isi = 11'h5;
                11'd197  : isi = 11'h5;
                11'd198  : isi = 11'h5;
                11'd199  : isi = 11'h5;
                11'd200  : isi = 11'h5;
                11'd201  : isi = 11'h5;
                11'd202  : isi = 11'h5;
                11'd203  : isi = 11'h5;
                11'd204  : isi = 11'h4;
                11'd205  : isi = 11'h4;
                11'd206  : isi = 11'h4;
                11'd207  : isi = 11'h4;
                11'd208  : isi = 11'h4;
                11'd209  : isi = 11'h4;
                11'd210  : isi = 11'h4;
                11'd211  : isi = 11'h4;
                11'd212  : isi = 11'h4;
                11'd213  : isi = 11'h4;
                11'd214  : isi = 11'h4;
                11'd215  : isi = 11'h4;
                11'd216  : isi = 11'h4;
                11'd217  : isi = 11'h4;
                11'd218  : isi = 11'h4;
                11'd219  : isi = 11'h4;
                11'd220  : isi = 11'h4;
                11'd221  : isi = 11'h4;
                11'd222  : isi = 11'h4;
                11'd223  : isi = 11'h4;
                11'd224  : isi = 11'h4;
                11'd225  : isi = 11'h4;
                11'd226  : isi = 11'h4;
                11'd227  : isi = 11'h4;
                11'd228  : isi = 11'h4;
                11'd229  : isi = 11'h4;
                11'd230  : isi = 11'h4;
                11'd231  : isi = 11'h4;
                11'd232  : isi = 11'h4;
                11'd233  : isi = 11'h4;
                11'd234  : isi = 11'h4;
                11'd235  : isi = 11'h4;
                11'd236  : isi = 11'h4;
                11'd237  : isi = 11'h4;
                11'd238  : isi = 11'h4;
                11'd239  : isi = 11'h4;
                11'd240  : isi = 11'h4;
                11'd241  : isi = 11'h4;
                11'd242  : isi = 11'h4;
                11'd243  : isi = 11'h4;
                11'd244  : isi = 11'h4;
                11'd245  : isi = 11'h4;
                11'd246  : isi = 11'h4;
                11'd247  : isi = 11'h4;
                11'd248  : isi = 11'h4;
                11'd249  : isi = 11'h4;
                11'd250  : isi = 11'h4;
                11'd251  : isi = 11'h4;
                11'd252  : isi = 11'h4;
                11'd253  : isi = 11'h4;
                11'd254  : isi = 11'h4;
                11'd255  : isi = 11'h4;
                11'd256  : isi = 11'h3;
                11'd257  : isi = 11'h3;
                11'd258  : isi = 11'h3;
                11'd259  : isi = 11'h3;
                11'd260  : isi = 11'h3;
                11'd261  : isi = 11'h3;
                11'd262  : isi = 11'h3;
                11'd263  : isi = 11'h3;
                11'd264  : isi = 11'h3;
                11'd265  : isi = 11'h3;
                11'd266  : isi = 11'h3;
                11'd267  : isi = 11'h3;
                11'd268  : isi = 11'h3;
                11'd269  : isi = 11'h3;
                11'd270  : isi = 11'h3;
                11'd271  : isi = 11'h3;
                11'd272  : isi = 11'h3;
                11'd273  : isi = 11'h3;
                11'd274  : isi = 11'h3;
                11'd275  : isi = 11'h3;
                11'd276  : isi = 11'h3;
                11'd277  : isi = 11'h3;
                11'd278  : isi = 11'h3;
                11'd279  : isi = 11'h3;
                11'd280  : isi = 11'h3;
                11'd281  : isi = 11'h3;
                11'd282  : isi = 11'h3;
                11'd283  : isi = 11'h3;
                11'd284  : isi = 11'h3;
                11'd285  : isi = 11'h3;
                11'd286  : isi = 11'h3;
                11'd287  : isi = 11'h3;
                11'd288  : isi = 11'h3;
                11'd289  : isi = 11'h3;
                11'd290  : isi = 11'h3;
                11'd291  : isi = 11'h3;
                11'd292  : isi = 11'h3;
                11'd293  : isi = 11'h3;
                11'd294  : isi = 11'h3;
                11'd295  : isi = 11'h3;
                11'd296  : isi = 11'h3;
                11'd297  : isi = 11'h3;
                11'd298  : isi = 11'h3;
                11'd299  : isi = 11'h3;
                11'd300  : isi = 11'h3;
                11'd301  : isi = 11'h3;
                11'd302  : isi = 11'h3;
                11'd303  : isi = 11'h3;
                11'd304  : isi = 11'h3;
                11'd305  : isi = 11'h3;
                11'd306  : isi = 11'h3;
                11'd307  : isi = 11'h3;
                11'd308  : isi = 11'h3;
                11'd309  : isi = 11'h3;
                11'd310  : isi = 11'h3;
                11'd311  : isi = 11'h3;
                11'd312  : isi = 11'h3;
                11'd313  : isi = 11'h3;
                11'd314  : isi = 11'h3;
                11'd315  : isi = 11'h3;
                11'd316  : isi = 11'h3;
                11'd317  : isi = 11'h3;
                11'd318  : isi = 11'h3;
                11'd319  : isi = 11'h3;
                11'd320  : isi = 11'h3;
                11'd321  : isi = 11'h3;
                11'd322  : isi = 11'h3;
                11'd323  : isi = 11'h3;
                11'd324  : isi = 11'h3;
                11'd325  : isi = 11'h3;
                11'd326  : isi = 11'h3;
                11'd327  : isi = 11'h3;
                11'd328  : isi = 11'h3;
                11'd329  : isi = 11'h3;
                11'd330  : isi = 11'h3;
                11'd331  : isi = 11'h3;
                11'd332  : isi = 11'h3;
                11'd333  : isi = 11'h3;
                11'd334  : isi = 11'h3;
                11'd335  : isi = 11'h3;
                11'd336  : isi = 11'h3;
                11'd337  : isi = 11'h3;
                11'd338  : isi = 11'h3;
                11'd339  : isi = 11'h3;
                11'd340  : isi = 11'h3;
                11'd341  : isi = 11'h2;
                11'd342  : isi = 11'h2;
                11'd343  : isi = 11'h2;
                11'd344  : isi = 11'h2;
                11'd345  : isi = 11'h2;
                11'd346  : isi = 11'h2;
                11'd347  : isi = 11'h2;
                11'd348  : isi = 11'h2;
                11'd349  : isi = 11'h2;
                11'd350  : isi = 11'h2;
                11'd351  : isi = 11'h2;
                11'd352  : isi = 11'h2;
                11'd353  : isi = 11'h2;
                11'd354  : isi = 11'h2;
                11'd355  : isi = 11'h2;
                11'd356  : isi = 11'h2;
                11'd357  : isi = 11'h2;
                11'd358  : isi = 11'h2;
                11'd359  : isi = 11'h2;
                11'd360  : isi = 11'h2;
                11'd361  : isi = 11'h2;
                11'd362  : isi = 11'h2;
                11'd363  : isi = 11'h2;
                11'd364  : isi = 11'h2;
                11'd365  : isi = 11'h2;
                11'd366  : isi = 11'h2;
                11'd367  : isi = 11'h2;
                11'd368  : isi = 11'h2;
                11'd369  : isi = 11'h2;
                11'd370  : isi = 11'h2;
                11'd371  : isi = 11'h2;
                11'd372  : isi = 11'h2;
                11'd373  : isi = 11'h2;
                11'd374  : isi = 11'h2;
                11'd375  : isi = 11'h2;
                11'd376  : isi = 11'h2;
                11'd377  : isi = 11'h2;
                11'd378  : isi = 11'h2;
                11'd379  : isi = 11'h2;
                11'd380  : isi = 11'h2;
                11'd381  : isi = 11'h2;
                11'd382  : isi = 11'h2;
                11'd383  : isi = 11'h2;
                11'd384  : isi = 11'h2;
                11'd385  : isi = 11'h2;
                11'd386  : isi = 11'h2;
                11'd387  : isi = 11'h2;
                11'd388  : isi = 11'h2;
                11'd389  : isi = 11'h2;
                11'd390  : isi = 11'h2;
                11'd391  : isi = 11'h2;
                11'd392  : isi = 11'h2;
                11'd393  : isi = 11'h2;
                11'd394  : isi = 11'h2;
                11'd395  : isi = 11'h2;
                11'd396  : isi = 11'h2;
                11'd397  : isi = 11'h2;
                11'd398  : isi = 11'h2;
                11'd399  : isi = 11'h2;
                11'd400  : isi = 11'h2;
                11'd401  : isi = 11'h2;
                11'd402  : isi = 11'h2;
                11'd403  : isi = 11'h2;
                11'd404  : isi = 11'h2;
                11'd405  : isi = 11'h2;
                11'd406  : isi = 11'h2;
                11'd407  : isi = 11'h2;
                11'd408  : isi = 11'h2;
                11'd409  : isi = 11'h2;
                11'd410  : isi = 11'h2;
                11'd411  : isi = 11'h2;
                11'd412  : isi = 11'h2;
                11'd413  : isi = 11'h2;
                11'd414  : isi = 11'h2;
                11'd415  : isi = 11'h2;
                11'd416  : isi = 11'h2;
                11'd417  : isi = 11'h2;
                11'd418  : isi = 11'h2;
                11'd419  : isi = 11'h2;
                11'd420  : isi = 11'h2;
                11'd421  : isi = 11'h2;
                11'd422  : isi = 11'h2;
                11'd423  : isi = 11'h2;
                11'd424  : isi = 11'h2;
                11'd425  : isi = 11'h2;
                11'd426  : isi = 11'h2;
                11'd427  : isi = 11'h2;
                11'd428  : isi = 11'h2;
                11'd429  : isi = 11'h2;
                11'd430  : isi = 11'h2;
                11'd431  : isi = 11'h2;
                11'd432  : isi = 11'h2;
                11'd433  : isi = 11'h2;
                11'd434  : isi = 11'h2;
                11'd435  : isi = 11'h2;
                11'd436  : isi = 11'h2;
                11'd437  : isi = 11'h2;
                11'd438  : isi = 11'h2;
                11'd439  : isi = 11'h2;
                11'd440  : isi = 11'h2;
                11'd441  : isi = 11'h2;
                11'd442  : isi = 11'h2;
                11'd443  : isi = 11'h2;
                11'd444  : isi = 11'h2;
                11'd445  : isi = 11'h2;
                11'd446  : isi = 11'h2;
                11'd447  : isi = 11'h2;
                11'd448  : isi = 11'h2;
                11'd449  : isi = 11'h2;
                11'd450  : isi = 11'h2;
                11'd451  : isi = 11'h2;
                11'd452  : isi = 11'h2;
                11'd453  : isi = 11'h2;
                11'd454  : isi = 11'h2;
                11'd455  : isi = 11'h2;
                11'd456  : isi = 11'h2;
                11'd457  : isi = 11'h2;
                11'd458  : isi = 11'h2;
                11'd459  : isi = 11'h2;
                11'd460  : isi = 11'h2;
                11'd461  : isi = 11'h2;
                11'd462  : isi = 11'h2;
                11'd463  : isi = 11'h2;
                11'd464  : isi = 11'h2;
                11'd465  : isi = 11'h2;
                11'd466  : isi = 11'h2;
                11'd467  : isi = 11'h2;
                11'd468  : isi = 11'h2;
                11'd469  : isi = 11'h2;
                11'd470  : isi = 11'h2;
                11'd471  : isi = 11'h2;
                11'd472  : isi = 11'h2;
                11'd473  : isi = 11'h2;
                11'd474  : isi = 11'h2;
                11'd475  : isi = 11'h2;
                11'd476  : isi = 11'h2;
                11'd477  : isi = 11'h2;
                11'd478  : isi = 11'h2;
                11'd479  : isi = 11'h2;
                11'd480  : isi = 11'h2;
                11'd481  : isi = 11'h2;
                11'd482  : isi = 11'h2;
                11'd483  : isi = 11'h2;
                11'd484  : isi = 11'h2;
                11'd485  : isi = 11'h2;
                11'd486  : isi = 11'h2;
                11'd487  : isi = 11'h2;
                11'd488  : isi = 11'h2;
                11'd489  : isi = 11'h2;
                11'd490  : isi = 11'h2;
                11'd491  : isi = 11'h2;
                11'd492  : isi = 11'h2;
                11'd493  : isi = 11'h2;
                11'd494  : isi = 11'h2;
                11'd495  : isi = 11'h2;
                11'd496  : isi = 11'h2;
                11'd497  : isi = 11'h2;
                11'd498  : isi = 11'h2;
                11'd499  : isi = 11'h2;
                11'd500  : isi = 11'h2;
                11'd501  : isi = 11'h2;
                11'd502  : isi = 11'h2;
                11'd503  : isi = 11'h2;
                11'd504  : isi = 11'h2;
                11'd505  : isi = 11'h2;
                11'd506  : isi = 11'h2;
                11'd507  : isi = 11'h2;
                11'd508  : isi = 11'h2;
                11'd509  : isi = 11'h2;
                11'd510  : isi = 11'h2;
                11'd511  : isi = 11'h2;
                11'd512  : isi = 11'h1;
                11'd513  : isi = 11'h1;
                11'd514  : isi = 11'h1;
                11'd515  : isi = 11'h1;
                11'd516  : isi = 11'h1;
                11'd517  : isi = 11'h1;
                11'd518  : isi = 11'h1;
                11'd519  : isi = 11'h1;
                11'd520  : isi = 11'h1;
                11'd521  : isi = 11'h1;
                11'd522  : isi = 11'h1;
                11'd523  : isi = 11'h1;
                11'd524  : isi = 11'h1;
                11'd525  : isi = 11'h1;
                11'd526  : isi = 11'h1;
                11'd527  : isi = 11'h1;
                11'd528  : isi = 11'h1;
                11'd529  : isi = 11'h1;
                11'd530  : isi = 11'h1;
                11'd531  : isi = 11'h1;
                11'd532  : isi = 11'h1;
                11'd533  : isi = 11'h1;
                11'd534  : isi = 11'h1;
                11'd535  : isi = 11'h1;
                11'd536  : isi = 11'h1;
                11'd537  : isi = 11'h1;
                11'd538  : isi = 11'h1;
                11'd539  : isi = 11'h1;
                11'd540  : isi = 11'h1;
                11'd541  : isi = 11'h1;
                11'd542  : isi = 11'h1;
                11'd543  : isi = 11'h1;
                11'd544  : isi = 11'h1;
                11'd545  : isi = 11'h1;
                11'd546  : isi = 11'h1;
                11'd547  : isi = 11'h1;
                11'd548  : isi = 11'h1;
                11'd549  : isi = 11'h1;
                11'd550  : isi = 11'h1;
                11'd551  : isi = 11'h1;
                11'd552  : isi = 11'h1;
                11'd553  : isi = 11'h1;
                11'd554  : isi = 11'h1;
                11'd555  : isi = 11'h1;
                11'd556  : isi = 11'h1;
                11'd557  : isi = 11'h1;
                11'd558  : isi = 11'h1;
                11'd559  : isi = 11'h1;
                11'd560  : isi = 11'h1;
                11'd561  : isi = 11'h1;
                11'd562  : isi = 11'h1;
                11'd563  : isi = 11'h1;
                11'd564  : isi = 11'h1;
                11'd565  : isi = 11'h1;
                11'd566  : isi = 11'h1;
                11'd567  : isi = 11'h1;
                11'd568  : isi = 11'h1;
                11'd569  : isi = 11'h1;
                11'd570  : isi = 11'h1;
                11'd571  : isi = 11'h1;
                11'd572  : isi = 11'h1;
                11'd573  : isi = 11'h1;
                11'd574  : isi = 11'h1;
                11'd575  : isi = 11'h1;
                11'd576  : isi = 11'h1;
                11'd577  : isi = 11'h1;
                11'd578  : isi = 11'h1;
                11'd579  : isi = 11'h1;
                11'd580  : isi = 11'h1;
                11'd581  : isi = 11'h1;
                11'd582  : isi = 11'h1;
                11'd583  : isi = 11'h1;
                11'd584  : isi = 11'h1;
                11'd585  : isi = 11'h1;
                11'd586  : isi = 11'h1;
                11'd587  : isi = 11'h1;
                11'd588  : isi = 11'h1;
                11'd589  : isi = 11'h1;
                11'd590  : isi = 11'h1;
                11'd591  : isi = 11'h1;
                11'd592  : isi = 11'h1;
                11'd593  : isi = 11'h1;
                11'd594  : isi = 11'h1;
                11'd595  : isi = 11'h1;
                11'd596  : isi = 11'h1;
                11'd597  : isi = 11'h1;
                11'd598  : isi = 11'h1;
                11'd599  : isi = 11'h1;
                11'd600  : isi = 11'h1;
                11'd601  : isi = 11'h1;
                11'd602  : isi = 11'h1;
                11'd603  : isi = 11'h1;
                11'd604  : isi = 11'h1;
                11'd605  : isi = 11'h1;
                11'd606  : isi = 11'h1;
                11'd607  : isi = 11'h1;
                11'd608  : isi = 11'h1;
                11'd609  : isi = 11'h1;
                11'd610  : isi = 11'h1;
                11'd611  : isi = 11'h1;
                11'd612  : isi = 11'h1;
                11'd613  : isi = 11'h1;
                11'd614  : isi = 11'h1;
                11'd615  : isi = 11'h1;
                11'd616  : isi = 11'h1;
                11'd617  : isi = 11'h1;
                11'd618  : isi = 11'h1;
                11'd619  : isi = 11'h1;
                11'd620  : isi = 11'h1;
                11'd621  : isi = 11'h1;
                11'd622  : isi = 11'h1;
                11'd623  : isi = 11'h1;
                11'd624  : isi = 11'h1;
                11'd625  : isi = 11'h1;
                11'd626  : isi = 11'h1;
                11'd627  : isi = 11'h1;
                11'd628  : isi = 11'h1;
                11'd629  : isi = 11'h1;
                11'd630  : isi = 11'h1;
                11'd631  : isi = 11'h1;
                11'd632  : isi = 11'h1;
                11'd633  : isi = 11'h1;
                11'd634  : isi = 11'h1;
                11'd635  : isi = 11'h1;
                11'd636  : isi = 11'h1;
                11'd637  : isi = 11'h1;
                11'd638  : isi = 11'h1;
                11'd639  : isi = 11'h1;
                11'd640  : isi = 11'h1;
                11'd641  : isi = 11'h1;
                11'd642  : isi = 11'h1;
                11'd643  : isi = 11'h1;
                11'd644  : isi = 11'h1;
                11'd645  : isi = 11'h1;
                11'd646  : isi = 11'h1;
                11'd647  : isi = 11'h1;
                11'd648  : isi = 11'h1;
                11'd649  : isi = 11'h1;
                11'd650  : isi = 11'h1;
                11'd651  : isi = 11'h1;
                11'd652  : isi = 11'h1;
                11'd653  : isi = 11'h1;
                11'd654  : isi = 11'h1;
                11'd655  : isi = 11'h1;
                11'd656  : isi = 11'h1;
                11'd657  : isi = 11'h1;
                11'd658  : isi = 11'h1;
                11'd659  : isi = 11'h1;
                11'd660  : isi = 11'h1;
                11'd661  : isi = 11'h1;
                11'd662  : isi = 11'h1;
                11'd663  : isi = 11'h1;
                11'd664  : isi = 11'h1;
                11'd665  : isi = 11'h1;
                11'd666  : isi = 11'h1;
                11'd667  : isi = 11'h1;
                11'd668  : isi = 11'h1;
                11'd669  : isi = 11'h1;
                11'd670  : isi = 11'h1;
                11'd671  : isi = 11'h1;
                11'd672  : isi = 11'h1;
                11'd673  : isi = 11'h1;
                11'd674  : isi = 11'h1;
                11'd675  : isi = 11'h1;
                11'd676  : isi = 11'h1;
                11'd677  : isi = 11'h1;
                11'd678  : isi = 11'h1;
                11'd679  : isi = 11'h1;
                11'd680  : isi = 11'h1;
                11'd681  : isi = 11'h1;
                11'd682  : isi = 11'h1;
                11'd683  : isi = 11'h1;
                11'd684  : isi = 11'h1;
                11'd685  : isi = 11'h1;
                11'd686  : isi = 11'h1;
                11'd687  : isi = 11'h1;
                11'd688  : isi = 11'h1;
                11'd689  : isi = 11'h1;
                11'd690  : isi = 11'h1;
                11'd691  : isi = 11'h1;
                11'd692  : isi = 11'h1;
                11'd693  : isi = 11'h1;
                11'd694  : isi = 11'h1;
                11'd695  : isi = 11'h1;
                11'd696  : isi = 11'h1;
                11'd697  : isi = 11'h1;
                11'd698  : isi = 11'h1;
                11'd699  : isi = 11'h1;
                11'd700  : isi = 11'h1;
                11'd701  : isi = 11'h1;
                11'd702  : isi = 11'h1;
                11'd703  : isi = 11'h1;
                11'd704  : isi = 11'h1;
                11'd705  : isi = 11'h1;
                11'd706  : isi = 11'h1;
                11'd707  : isi = 11'h1;
                11'd708  : isi = 11'h1;
                11'd709  : isi = 11'h1;
                11'd710  : isi = 11'h1;
                11'd711  : isi = 11'h1;
                11'd712  : isi = 11'h1;
                11'd713  : isi = 11'h1;
                11'd714  : isi = 11'h1;
                11'd715  : isi = 11'h1;
                11'd716  : isi = 11'h1;
                11'd717  : isi = 11'h1;
                11'd718  : isi = 11'h1;
                11'd719  : isi = 11'h1;
                11'd720  : isi = 11'h1;
                11'd721  : isi = 11'h1;
                11'd722  : isi = 11'h1;
                11'd723  : isi = 11'h1;
                11'd724  : isi = 11'h1;
                11'd725  : isi = 11'h1;
                11'd726  : isi = 11'h1;
                11'd727  : isi = 11'h1;
                11'd728  : isi = 11'h1;
                11'd729  : isi = 11'h1;
                11'd730  : isi = 11'h1;
                11'd731  : isi = 11'h1;
                11'd732  : isi = 11'h1;
                11'd733  : isi = 11'h1;
                11'd734  : isi = 11'h1;
                11'd735  : isi = 11'h1;
                11'd736  : isi = 11'h1;
                11'd737  : isi = 11'h1;
                11'd738  : isi = 11'h1;
                11'd739  : isi = 11'h1;
                11'd740  : isi = 11'h1;
                11'd741  : isi = 11'h1;
                11'd742  : isi = 11'h1;
                11'd743  : isi = 11'h1;
                11'd744  : isi = 11'h1;
                11'd745  : isi = 11'h1;
                11'd746  : isi = 11'h1;
                11'd747  : isi = 11'h1;
                11'd748  : isi = 11'h1;
                11'd749  : isi = 11'h1;
                11'd750  : isi = 11'h1;
                11'd751  : isi = 11'h1;
                11'd752  : isi = 11'h1;
                11'd753  : isi = 11'h1;
                11'd754  : isi = 11'h1;
                11'd755  : isi = 11'h1;
                11'd756  : isi = 11'h1;
                11'd757  : isi = 11'h1;
                11'd758  : isi = 11'h1;
                11'd759  : isi = 11'h1;
                11'd760  : isi = 11'h1;
                11'd761  : isi = 11'h1;
                11'd762  : isi = 11'h1;
                11'd763  : isi = 11'h1;
                11'd764  : isi = 11'h1;
                11'd765  : isi = 11'h1;
                11'd766  : isi = 11'h1;
                11'd767  : isi = 11'h1;
                11'd768  : isi = 11'h1;
                11'd769  : isi = 11'h1;
                11'd770  : isi = 11'h1;
                11'd771  : isi = 11'h1;
                11'd772  : isi = 11'h1;
                11'd773  : isi = 11'h1;
                11'd774  : isi = 11'h1;
                11'd775  : isi = 11'h1;
                11'd776  : isi = 11'h1;
                11'd777  : isi = 11'h1;
                11'd778  : isi = 11'h1;
                11'd779  : isi = 11'h1;
                11'd780  : isi = 11'h1;
                11'd781  : isi = 11'h1;
                11'd782  : isi = 11'h1;
                11'd783  : isi = 11'h1;
                11'd784  : isi = 11'h1;
                11'd785  : isi = 11'h1;
                11'd786  : isi = 11'h1;
                11'd787  : isi = 11'h1;
                11'd788  : isi = 11'h1;
                11'd789  : isi = 11'h1;
                11'd790  : isi = 11'h1;
                11'd791  : isi = 11'h1;
                11'd792  : isi = 11'h1;
                11'd793  : isi = 11'h1;
                11'd794  : isi = 11'h1;
                11'd795  : isi = 11'h1;
                11'd796  : isi = 11'h1;
                11'd797  : isi = 11'h1;
                11'd798  : isi = 11'h1;
                11'd799  : isi = 11'h1;
                11'd800  : isi = 11'h1;
                11'd801  : isi = 11'h1;
                11'd802  : isi = 11'h1;
                11'd803  : isi = 11'h1;
                11'd804  : isi = 11'h1;
                11'd805  : isi = 11'h1;
                11'd806  : isi = 11'h1;
                11'd807  : isi = 11'h1;
                11'd808  : isi = 11'h1;
                11'd809  : isi = 11'h1;
                11'd810  : isi = 11'h1;
                11'd811  : isi = 11'h1;
                11'd812  : isi = 11'h1;
                11'd813  : isi = 11'h1;
                11'd814  : isi = 11'h1;
                11'd815  : isi = 11'h1;
                11'd816  : isi = 11'h1;
                11'd817  : isi = 11'h1;
                11'd818  : isi = 11'h1;
                11'd819  : isi = 11'h1;
                11'd820  : isi = 11'h1;
                11'd821  : isi = 11'h1;
                11'd822  : isi = 11'h1;
                11'd823  : isi = 11'h1;
                11'd824  : isi = 11'h1;
                11'd825  : isi = 11'h1;
                11'd826  : isi = 11'h1;
                11'd827  : isi = 11'h1;
                11'd828  : isi = 11'h1;
                11'd829  : isi = 11'h1;
                11'd830  : isi = 11'h1;
                11'd831  : isi = 11'h1;
                11'd832  : isi = 11'h1;
                11'd833  : isi = 11'h1;
                11'd834  : isi = 11'h1;
                11'd835  : isi = 11'h1;
                11'd836  : isi = 11'h1;
                11'd837  : isi = 11'h1;
                11'd838  : isi = 11'h1;
                11'd839  : isi = 11'h1;
                11'd840  : isi = 11'h1;
                11'd841  : isi = 11'h1;
                11'd842  : isi = 11'h1;
                11'd843  : isi = 11'h1;
                11'd844  : isi = 11'h1;
                11'd845  : isi = 11'h1;
                11'd846  : isi = 11'h1;
                11'd847  : isi = 11'h1;
                11'd848  : isi = 11'h1;
                11'd849  : isi = 11'h1;
                11'd850  : isi = 11'h1;
                11'd851  : isi = 11'h1;
                11'd852  : isi = 11'h1;
                11'd853  : isi = 11'h1;
                11'd854  : isi = 11'h1;
                11'd855  : isi = 11'h1;
                11'd856  : isi = 11'h1;
                11'd857  : isi = 11'h1;
                11'd858  : isi = 11'h1;
                11'd859  : isi = 11'h1;
                11'd860  : isi = 11'h1;
                11'd861  : isi = 11'h1;
                11'd862  : isi = 11'h1;
                11'd863  : isi = 11'h1;
                11'd864  : isi = 11'h1;
                11'd865  : isi = 11'h1;
                11'd866  : isi = 11'h1;
                11'd867  : isi = 11'h1;
                11'd868  : isi = 11'h1;
                11'd869  : isi = 11'h1;
                11'd870  : isi = 11'h1;
                11'd871  : isi = 11'h1;
                11'd872  : isi = 11'h1;
                11'd873  : isi = 11'h1;
                11'd874  : isi = 11'h1;
                11'd875  : isi = 11'h1;
                11'd876  : isi = 11'h1;
                11'd877  : isi = 11'h1;
                11'd878  : isi = 11'h1;
                11'd879  : isi = 11'h1;
                11'd880  : isi = 11'h1;
                11'd881  : isi = 11'h1;
                11'd882  : isi = 11'h1;
                11'd883  : isi = 11'h1;
                11'd884  : isi = 11'h1;
                11'd885  : isi = 11'h1;
                11'd886  : isi = 11'h1;
                11'd887  : isi = 11'h1;
                11'd888  : isi = 11'h1;
                11'd889  : isi = 11'h1;
                11'd890  : isi = 11'h1;
                11'd891  : isi = 11'h1;
                11'd892  : isi = 11'h1;
                11'd893  : isi = 11'h1;
                11'd894  : isi = 11'h1;
                11'd895  : isi = 11'h1;
                11'd896  : isi = 11'h1;
                11'd897  : isi = 11'h1;
                11'd898  : isi = 11'h1;
                11'd899  : isi = 11'h1;
                11'd900  : isi = 11'h1;
                11'd901  : isi = 11'h1;
                11'd902  : isi = 11'h1;
                11'd903  : isi = 11'h1;
                11'd904  : isi = 11'h1;
                11'd905  : isi = 11'h1;
                11'd906  : isi = 11'h1;
                11'd907  : isi = 11'h1;
                11'd908  : isi = 11'h1;
                11'd909  : isi = 11'h1;
                11'd910  : isi = 11'h1;
                11'd911  : isi = 11'h1;
                11'd912  : isi = 11'h1;
                11'd913  : isi = 11'h1;
                11'd914  : isi = 11'h1;
                11'd915  : isi = 11'h1;
                11'd916  : isi = 11'h1;
                11'd917  : isi = 11'h1;
                11'd918  : isi = 11'h1;
                11'd919  : isi = 11'h1;
                11'd920  : isi = 11'h1;
                11'd921  : isi = 11'h1;
                11'd922  : isi = 11'h1;
                11'd923  : isi = 11'h1;
                11'd924  : isi = 11'h1;
                11'd925  : isi = 11'h1;
                11'd926  : isi = 11'h1;
                11'd927  : isi = 11'h1;
                11'd928  : isi = 11'h1;
                11'd929  : isi = 11'h1;
                11'd930  : isi = 11'h1;
                11'd931  : isi = 11'h1;
                11'd932  : isi = 11'h1;
                11'd933  : isi = 11'h1;
                11'd934  : isi = 11'h1;
                11'd935  : isi = 11'h1;
                11'd936  : isi = 11'h1;
                11'd937  : isi = 11'h1;
                11'd938  : isi = 11'h1;
                11'd939  : isi = 11'h1;
                11'd940  : isi = 11'h1;
                11'd941  : isi = 11'h1;
                11'd942  : isi = 11'h1;
                11'd943  : isi = 11'h1;
                11'd944  : isi = 11'h1;
                11'd945  : isi = 11'h1;
                11'd946  : isi = 11'h1;
                11'd947  : isi = 11'h1;
                11'd948  : isi = 11'h1;
                11'd949  : isi = 11'h1;
                11'd950  : isi = 11'h1;
                11'd951  : isi = 11'h1;
                11'd952  : isi = 11'h1;
                11'd953  : isi = 11'h1;
                11'd954  : isi = 11'h1;
                11'd955  : isi = 11'h1;
                11'd956  : isi = 11'h1;
                11'd957  : isi = 11'h1;
                11'd958  : isi = 11'h1;
                11'd959  : isi = 11'h1;
                11'd960  : isi = 11'h1;
                11'd961  : isi = 11'h1;
                11'd962  : isi = 11'h1;
                11'd963  : isi = 11'h1;
                11'd964  : isi = 11'h1;
                11'd965  : isi = 11'h1;
                11'd966  : isi = 11'h1;
                11'd967  : isi = 11'h1;
                11'd968  : isi = 11'h1;
                11'd969  : isi = 11'h1;
                11'd970  : isi = 11'h1;
                11'd971  : isi = 11'h1;
                11'd972  : isi = 11'h1;
                11'd973  : isi = 11'h1;
                11'd974  : isi = 11'h1;
                11'd975  : isi = 11'h1;
                11'd976  : isi = 11'h1;
                11'd977  : isi = 11'h1;
                11'd978  : isi = 11'h1;
                11'd979  : isi = 11'h1;
                11'd980  : isi = 11'h1;
                11'd981  : isi = 11'h1;
                11'd982  : isi = 11'h1;
                11'd983  : isi = 11'h1;
                11'd984  : isi = 11'h1;
                11'd985  : isi = 11'h1;
                11'd986  : isi = 11'h1;
                11'd987  : isi = 11'h1;
                11'd988  : isi = 11'h1;
                11'd989  : isi = 11'h1;
                11'd990  : isi = 11'h1;
                11'd991  : isi = 11'h1;
                11'd992  : isi = 11'h1;
                11'd993  : isi = 11'h1;
                11'd994  : isi = 11'h1;
                11'd995  : isi = 11'h1;
                11'd996  : isi = 11'h1;
                11'd997  : isi = 11'h1;
                11'd998  : isi = 11'h1;
                11'd999  : isi = 11'h1;
                11'd1000  : isi = 11'h1;
                11'd1001  : isi = 11'h1;
                11'd1002  : isi = 11'h1;
                11'd1003  : isi = 11'h1;
                11'd1004  : isi = 11'h1;
                11'd1005  : isi = 11'h1;
                11'd1006  : isi = 11'h1;
                11'd1007  : isi = 11'h1;
                11'd1008  : isi = 11'h1;
                11'd1009  : isi = 11'h1;
                11'd1010  : isi = 11'h1;
                11'd1011  : isi = 11'h1;
                11'd1012  : isi = 11'h1;
                11'd1013  : isi = 11'h1;
                11'd1014  : isi = 11'h1;
                11'd1015  : isi = 11'h1;
                11'd1016  : isi = 11'h1;
                11'd1017  : isi = 11'h1;
                11'd1018  : isi = 11'h1;
                11'd1019  : isi = 11'h1;
                11'd1020  : isi = 11'h1;
                11'd1021  : isi = 11'h1;
                11'd1022  : isi = 11'h1;
                11'd1023  : isi = 11'h1;
    endcase
    end

			
endmodule
